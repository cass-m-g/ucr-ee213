V1 1 0 15
R1 1 2 2.7K
R2 2 0 5k
R35 2 3 1MEG
RZ 3 0 10k
.end
