* Test netlist 2 -- voltage devider

R1 1 2 1000 
R2 2 0 1000
Vs1 1 0 2

.end
