R1 1 0 5
G2 1 0 1 2 2
R3 1 2 6
R4 2 0 8
Is 0 2 PWL(0 0 
+ 17ns 1 
+ 32ns 2
+ 47ns 3
+ 62ns 4
+ 77ns 5
+ 92ns 6
+ 107ns 7
+ 122ns 8
+ 137ns 9
+ 152ns 10
+ )


.end
