R1 N1 N2 1.0
R2 N2 N3 1.0
R3 N1 N2 1.0
C1_0 N1_0 0 1.15e-12
.end